/*
 *  EV3_mruby_common.cdl
 *  
 */

import(<kernel.cdl>);

/* mrubyの本体 */
import(<tMruby.cdl>);

import(<tUltrasonicSensor.cdl>);
import(<tColorSensor.cdl>);
import(<tTouchSensor.cdl>);
import(<tGyroSensor.cdl>);

import(<tMotor.cdl>);

import(<tLCD.cdl>);
import(<tLED.cdl>);
import(<tButton.cdl>);
import(<tBattery.cdl>);
import(<tSpeaker.cdl>);

import(<tEV3Platform.cdl>);
import(<tBalancer.cdl>);

import("tReset.cdl");

/*
 * シグニチャプラグイン MrubyBridgePlugin の呼び出し。
 */
generate( MrubyBridgePlugin, sKernel, "" );

generate( MrubyBridgePlugin, sMotor, "" );

generate( MrubyBridgePlugin, sLCD, "" );
generate( MrubyBridgePlugin, sLED, "" );
generate( MrubyBridgePlugin, sButton, "" );
generate( MrubyBridgePlugin, sBattery, "" );
generate( MrubyBridgePlugin, sSpeaker, "" );

generate( MrubyBridgePlugin, sUltrasonicSensor, "" );
generate( MrubyBridgePlugin, sGyroSensor, "" );
generate( MrubyBridgePlugin, sColorSensor, "" );
generate( MrubyBridgePlugin, sTouchSensor, "" );

generate( MrubyBridgePlugin, sBalancer, "" );

[domain(HRP2, "trusted")]
region rDomainEV3{
	//Kernel
	cell tKernel HRP2Kernel{
	};
    //Motor
	cell tMotor MotorA{
		port = C_EXP("EV3_PORT_A");
	};
	cell tMotor MotorB{
		port = C_EXP("EV3_PORT_B");
	};
	cell tMotor MotorC{
		port = C_EXP("EV3_PORT_C");
	};
	cell tMotor MotorD{
		port = C_EXP("EV3_PORT_D");
	};
	//LCD
	cell tLCD LCD{
		cButton = Button.eButton;
	};
	//LED
	cell tLED LED{
	};
	//Button
	cell tButton Button{
	};
	//Battery
	cell tBattery Battery{
	};
	//Speaker
	cell tSpeaker Speaker{
	};
	//UltrasonicSensor
	cell tUltrasonicSensor UltrasonicSensor1{
		port = C_EXP("EV3_PORT_1");
	};
	cell tUltrasonicSensor UltrasonicSensor2{
		port = C_EXP("EV3_PORT_2");
	};
	cell tUltrasonicSensor UltrasonicSensor3{
		port = C_EXP("EV3_PORT_3");
	};
	cell tUltrasonicSensor UltrasonicSensor4{
		port = C_EXP("EV3_PORT_4");
	};
	//GyroSensor
	cell tGyroSensor GyroSensor1{
		port = C_EXP("EV3_PORT_1");
	};
	cell tGyroSensor GyroSensor2{
		port = C_EXP("EV3_PORT_2");
	};
	cell tGyroSensor GyroSensor3{
		port = C_EXP("EV3_PORT_3");
	};
	cell tGyroSensor GyroSensor4{
		port = C_EXP("EV3_PORT_4");
	};
	//ColorSensor
	cell tColorSensor ColorSensor1{
		port = C_EXP("EV3_PORT_1");
	};
	cell tColorSensor ColorSensor2{
		port = C_EXP("EV3_PORT_2");
	};
	cell tColorSensor ColorSensor3{
		port = C_EXP("EV3_PORT_3");
	};
	cell tColorSensor ColorSensor4{
		port = C_EXP("EV3_PORT_4");
	};
	//TouchSensor
	cell tTouchSensor TouchSensor1{
		port = C_EXP("EV3_PORT_1");
	};
	cell tTouchSensor TouchSensor2{
		port = C_EXP("EV3_PORT_2");
	};
	cell tTouchSensor TouchSensor3{
		port = C_EXP("EV3_PORT_3");
	};
	cell tTouchSensor TouchSensor4{
		port = C_EXP("EV3_PORT_4");
	};
	
	cell tBalancer Balancer{
		
	};

};
