/*
 *  tEV3Sample.cdl
 *
 */

import("VM1.cdl");
