/*
 *   TOPPERS Software
 *       Toyohashi Open Platform for Embedded Real-Time Systems
 *
 *   Copyright (C) 2010-2011 by Embedded and Real-Time Systems Laboratory
 *               Graduate School of Information Science, Nagoya Univ., JAPAN
 *
 *   �嵭����Ԥϡ��ʲ���(1)��(4)�ξ������������˸¤ꡤ�ܥ��եȥ���
 *   �����ܥ��եȥ���������Ѥ�����Τ�ޤࡥ�ʲ�Ʊ���ˤ���ѡ�ʣ������
 *   �ѡ������ۡʰʲ������ѤȸƤ֡ˤ��뤳�Ȥ�̵���ǵ������롥
 *   (1) �ܥ��եȥ������򥽡��������ɤη������Ѥ�����ˤϡ��嵭������
 *       ��ɽ�����������Ѿ�浪��Ӳ�����̵�ݾڵ��꤬�����Τޤޤη��ǥ���
 *       ����������˴ޤޤ�Ƥ��뤳�ȡ�
 *   (2) �ܥ��եȥ������򡤥饤�֥������ʤɡ�¾�Υ��եȥ�������ȯ�˻�
 *       �ѤǤ�����Ǻ����ۤ�����ˤϡ������ۤ�ȼ���ɥ�����ȡ�����
 *       �ԥޥ˥奢��ʤɡˤˡ��嵭�����ɽ�����������Ѿ�浪��Ӳ���
 *       ��̵�ݾڵ����Ǻܤ��뤳�ȡ�
 *   (3) �ܥ��եȥ������򡤵�����Ȥ߹���ʤɡ�¾�Υ��եȥ�������ȯ�˻�
 *       �ѤǤ��ʤ����Ǻ����ۤ�����ˤϡ����Τ����줫�ξ�����������
 *       �ȡ�
 *     (a) �����ۤ�ȼ���ɥ�����ȡ����Ѽԥޥ˥奢��ʤɡˤˡ��嵭����
 *         �ɽ�����������Ѿ�浪��Ӳ�����̵�ݾڵ����Ǻܤ��뤳�ȡ�
 *     (b) �����ۤη��֤��̤�������ˡ�ˤ�äơ�TOPPERS�ץ������Ȥ�
 *         ��𤹤뤳�ȡ�
 *   (4) �ܥ��եȥ����������Ѥˤ��ľ��Ū�ޤ��ϴ���Ū�������뤤���ʤ�»
 *       ������⡤�嵭����Ԥ����TOPPERS�ץ������Ȥ����դ��뤳�ȡ�
 *       �ޤ����ܥ��եȥ������Υ桼���ޤ��ϥ���ɥ桼������Τ����ʤ���
 *       ͳ�˴�Ť����ᤫ��⡤�嵭����Ԥ����TOPPERS�ץ������Ȥ�
 *       ���դ��뤳�ȡ�
 *
 *   �ܥ��եȥ������ϡ�̵�ݾڤ��󶡤���Ƥ����ΤǤ��롥�嵭����Ԥ�
 *   ���TOPPERS�ץ������Ȥϡ��ܥ��եȥ������˴ؤ��ơ�����λ�����Ū
 *   ���Ф���Ŭ������ޤ�ơ������ʤ��ݾڤ�Ԥ�ʤ����ޤ����ܥ��եȥ���
 *   �������Ѥˤ��ľ��Ū�ޤ��ϴ���Ū�������������ʤ�»���˴ؤ��Ƥ⡤��
 *   ����Ǥ�����ʤ���
 *
 */

/*
 *  ��Ω����׻��Τ���Υ����˥���
 */
signature sBalancer {
	/* ��Ω����Τ���Υѥ�᡼����׻����� */
	/*void control([in] int16_t forward, [in] int16_t turn,
                 [in] uint16_t gyro, [in] uint16_t gyroOffset,
                 [in] int32_t leftRevolution, [in] int32_t rightRevolution,
                 [in] uint16_t battery,
                 [out] int8_t *pwm_l, [out] int8_t *pwm_r);*/
	void control([in] float32_t forward, [in] float32_t turn,
                 [in] float32_t gyro, [in] float32_t gyroOffset,
                 [in] float32_t leftRevolution, [in] float32_t rightRevolution,
                 [in] float32_t battery,
                 [out] int8_t *pwm_l, [out] int8_t *pwm_r);
	void init(void);
};

/*
 *  �Х�󥵤����
 */
[singleton]
celltype tBalancer{
	entry sBalancer eBalancer;
//    [inline] entry sBalancer eBalancer;
//    [inline] entry sInitializeRoutineBody eInitialize;

    FACTORY {
        /* ��Ω����׻��Τ���Υ饤�֥�����ɥ⥸�塼��˴ޤ�� */
//       write("$ct$_tecsgen.h", "#include \"balancer.h\"");
        write("Makefile.tecsgen", "SYSSVC_COBJS := balancer.o balancer_param.o $(SYSSVC_COBJS)");
//        write("Makefile.tecsgen", "SYSSVC_COBJS :=  balancer_param.o $(SYSSVC_COBJS)");
        write("Makefile.tecsgen", "INCLUDES := -I$(SRCDIR)/tecs_lib/mindstorms_ev3/balancer $(INCLUDES)");
        write("Makefile.tecsgen", "vpath %.c $(SRCDIR)/tecs_lib/mindstorms_ev3/balancer");
	write("tecsgen.cfg","ATT\_MOD\(\"balancer.o\"\);");
	write("tecsgen.cfg","ATT\_MOD\(\"balancer_param.o\"\);");
    };
};
